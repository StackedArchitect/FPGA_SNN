// Automatically generated weight parameters for CONV_BIAS
// Bit width: 8
// Generated from quantize_weights.py

// Total weights: 4
// Original shape: (4,)

parameter [7:0] CONV_BIAS [0:3] = '{
    8'h02, 8'hF6, 8'h00, 8'hF6
};

