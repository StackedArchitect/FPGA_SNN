// Automatically generated weight parameters for FC_WEIGHTS
// Bit width: 8
// Generated from quantize_weights.py

// Total weights: 6760
// Original shape: (10, 676)

parameter [7:0] FC_WEIGHTS [0:6759] = '{
    8'h00, 8'h01, 8'h01, 8'h00, 8'h01, 8'h01, 8'h02, 8'h01,
    8'h02, 8'h01, 8'h01, 8'h00, 8'h01, 8'h01, 8'h01, 8'h01,
    8'h02, 8'h02, 8'h02, 8'h02, 8'h01, 8'h03, 8'h01, 8'h01,
    8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h00, 8'hFF,
    8'h01, 8'h01, 8'hFD, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h01,
    8'h01, 8'h00, 8'h00, 8'hFE, 8'h00, 8'hFF, 8'hFD, 8'hFB,
    8'hFA, 8'hFB, 8'hFF, 8'h01, 8'h01, 8'h01, 8'h00, 8'hFF,
    8'h00, 8'hFF, 8'hFE, 8'hFD, 8'hFA, 8'hF9, 8'hFB, 8'hFE,
    8'h01, 8'h01, 8'h02, 8'hFF, 8'h01, 8'h01, 8'hFD, 8'h01,
    8'h02, 8'hFD, 8'hFA, 8'hFA, 8'hFD, 8'h00, 8'h00, 8'h02,
    8'hFE, 8'hFF, 8'hFD, 8'hFE, 8'h00, 8'h02, 8'h00, 8'h00,
    8'hFF, 8'hFE, 8'h00, 8'h01, 8'h00, 8'hFF, 8'hFC, 8'hFE,
    8'hFF, 8'h01, 8'h02, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00,
    8'h01, 8'h00, 8'h00, 8'hFB, 8'hFB, 8'h00, 8'h02, 8'h04,
    8'h04, 8'h02, 8'h01, 8'h01, 8'h00, 8'h02, 8'h00, 8'hFF,
    8'hFE, 8'hFB, 8'hFE, 8'h06, 8'h05, 8'h04, 8'h01, 8'h01,
    8'h01, 8'h02, 8'h01, 8'h01, 8'h00, 8'hFF, 8'hFC, 8'hFF,
    8'h01, 8'h02, 8'h02, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01,
    8'h01, 8'h01, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h01,
    8'h01, 8'h01, 8'h00, 8'h00, 8'h01, 8'h00, 8'h01, 8'h01,
    8'h00, 8'hFF, 8'h01, 8'h01, 8'h01, 8'h00, 8'h00, 8'h00,
    8'h01, 8'hFF, 8'h00, 8'hFF, 8'hFD, 8'hFA, 8'hFE, 8'hFF,
    8'hFA, 8'hFB, 8'hFE, 8'hFE, 8'hFE, 8'h02, 8'hFE, 8'hFE,
    8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFE, 8'hFE, 8'hFF,
    8'hFF, 8'h00, 8'hFE, 8'h01, 8'hFC, 8'h01, 8'h01, 8'h01,
    8'hFF, 8'h00, 8'hFF, 8'h00, 8'h00, 8'h00, 8'hFE, 8'hFC,
    8'hFE, 8'hFF, 8'h02, 8'hFF, 8'h00, 8'hFF, 8'h01, 8'h01,
    8'h01, 8'hFF, 8'hFF, 8'h00, 8'hFA, 8'h03, 8'hFF, 8'h01,
    8'h01, 8'h02, 8'h00, 8'h01, 8'h00, 8'hFF, 8'h00, 8'hFF,
    8'h01, 8'hFD, 8'h02, 8'hFF, 8'h01, 8'h01, 8'h01, 8'h01,
    8'h00, 8'hFF, 8'hFF, 8'h01, 8'h01, 8'h01, 8'hFE, 8'h02,
    8'hFF, 8'h03, 8'h03, 8'h03, 8'h01, 8'hFE, 8'hFC, 8'h00,
    8'h00, 8'h02, 8'h02, 8'hFF, 8'hFE, 8'h00, 8'h01, 8'h02,
    8'h03, 8'h00, 8'hFA, 8'hFD, 8'h00, 8'h01, 8'h02, 8'h03,
    8'hFE, 8'h00, 8'h01, 8'h01, 8'h01, 8'h01, 8'h00, 8'hFD,
    8'hFE, 8'hFF, 8'h00, 8'h01, 8'h02, 8'hFF, 8'hFB, 8'h01,
    8'hFF, 8'h01, 8'h01, 8'h01, 8'hFF, 8'h00, 8'h00, 8'h00,
    8'h01, 8'h01, 8'hFB, 8'hFD, 8'hFF, 8'hFF, 8'h00, 8'h00,
    8'h00, 8'hFE, 8'h00, 8'hFF, 8'hFE, 8'h02, 8'h01, 8'h01,
    8'hFE, 8'hFB, 8'h02, 8'hFF, 8'hFF, 8'h00, 8'hFF, 8'h00,
    8'hFF, 8'hFE, 8'h00, 8'hFA, 8'h00, 8'hFD, 8'h02, 8'hFD,
    8'hFD, 8'hF9, 8'hFB, 8'hFB, 8'hF6, 8'hF9, 8'hF8, 8'hFC,
    8'hFD, 8'h00, 8'h03, 8'hFF, 8'hFC, 8'hFC, 8'hFF, 8'h00,
    8'hFF, 8'hFE, 8'hFE, 8'hFD, 8'hFE, 8'hFF, 8'hFF, 8'h02,
    8'hFC, 8'hFF, 8'h01, 8'h00, 8'hFF, 8'h00, 8'h00, 8'h00,
    8'h01, 8'hFF, 8'h00, 8'hFC, 8'hFF, 8'hFE, 8'h01, 8'h00,
    8'h00, 8'h00, 8'h00, 8'h02, 8'h00, 8'hFF, 8'h00, 8'h02,
    8'h00, 8'h04, 8'hFF, 8'h00, 8'h01, 8'hFF, 8'hFF, 8'h00,
    8'h01, 8'h03, 8'h01, 8'h00, 8'hFF, 8'hFD, 8'h04, 8'h01,
    8'h01, 8'h00, 8'hFE, 8'hFF, 8'hFE, 8'hFD, 8'hFF, 8'hFE,
    8'h02, 8'h01, 8'hFD, 8'h02, 8'h01, 8'h01, 8'h02, 8'h02,
    8'h00, 8'hFE, 8'hFD, 8'hFC, 8'h00, 8'hFF, 8'h02, 8'hFF,
    8'h00, 8'h01, 8'h02, 8'h01, 8'h03, 8'hFF, 8'hFC, 8'hFF,
    8'hFE, 8'h00, 8'h01, 8'hFF, 8'h00, 8'hFD, 8'h02, 8'h02,
    8'h00, 8'h00, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFE, 8'h00,
    8'hFF, 8'hFC, 8'hFD, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF,
    8'h01, 8'h00, 8'h01, 8'h02, 8'hFF, 8'hFC, 8'hFA, 8'hFD,
    8'h00, 8'h00, 8'hFF, 8'h01, 8'h00, 8'h03, 8'h03, 8'h02,
    8'h01, 8'h01, 8'hFF, 8'hFE, 8'h01, 8'hFF, 8'hFE, 8'hFD,
    8'h00, 8'h01, 8'h02, 8'h01, 8'h00, 8'h02, 8'h00, 8'hFF,
    8'h04, 8'hFD, 8'h01, 8'h00, 8'hFE, 8'h02, 8'h00, 8'h00,
    8'h02, 8'h00, 8'h01, 8'hF7, 8'hFD, 8'h02, 8'h01, 8'h00,
    8'hFD, 8'hFB, 8'hFB, 8'hFC, 8'hF6, 8'hF4, 8'hF7, 8'hF9,
    8'hFC, 8'h00, 8'h02, 8'h01, 8'h00, 8'h00, 8'hFD, 8'h02,
    8'h01, 8'h00, 8'h01, 8'h00, 8'hFC, 8'hFC, 8'hFF, 8'h00,
    8'h00, 8'hFF, 8'h01, 8'hFF, 8'hFE, 8'hFD, 8'hFE, 8'h01,
    8'h01, 8'h02, 8'hFD, 8'h01, 8'h02, 8'hFC, 8'hFB, 8'hFC,
    8'hFD, 8'hFB, 8'hFC, 8'hFF, 8'h00, 8'h00, 8'h02, 8'h01,
    8'hFC, 8'hF8, 8'h00, 8'h02, 8'hFF, 8'hFD, 8'hFC, 8'h00,
    8'h01, 8'h01, 8'h04, 8'h02, 8'h04, 8'h01, 8'hFD, 8'h03,
    8'hFD, 8'hFC, 8'hFE, 8'hFF, 8'hFF, 8'h00, 8'h02, 8'h01,
    8'h02, 8'h02, 8'hFF, 8'hF9, 8'h03, 8'hFE, 8'hFC, 8'hFB,
    8'hFD, 8'hFE, 8'h00, 8'h01, 8'hFF, 8'h00, 8'h02, 8'h00,
    8'hF5, 8'h01, 8'hFF, 8'hFE, 8'hFA, 8'hFE, 8'hFD, 8'hFD,
    8'hFE, 8'h00, 8'hFF, 8'h00, 8'hFE, 8'hFA, 8'hFB, 8'hFF,
    8'hFF, 8'hFD, 8'hFC, 8'hFE, 8'hFB, 8'hFA, 8'hFD, 8'hFF,
    8'hFE, 8'hFF, 8'h00, 8'hFE, 8'hFF, 8'hFF, 8'h00, 8'h00,
    8'hFB, 8'hFB, 8'hFD, 8'hFE, 8'hFE, 8'hFF, 8'h00, 8'hFD,
    8'hFC, 8'h00, 8'hFE, 8'hFE, 8'h02, 8'h00, 8'hFF, 8'hFF,
    8'hFD, 8'hFE, 8'h00, 8'hFE, 8'hFD, 8'h00, 8'h00, 8'h00,
    8'hFF, 8'h02, 8'h03, 8'h01, 8'hFF, 8'hFE, 8'hFE, 8'hFE,
    8'hFC, 8'h03, 8'hFB, 8'hFE, 8'h02, 8'h02, 8'h02, 8'h03,
    8'h02, 8'h01, 8'hFF, 8'hFE, 8'h01, 8'hFC, 8'hFC, 8'hFD,
    8'h01, 8'hFF, 8'h00, 8'hFE, 8'h00, 8'h00, 8'hFF, 8'hFE,
    8'hFA, 8'hFA, 8'hFB, 8'hFB, 8'h02, 8'h02, 8'h01, 8'h02,
    8'h02, 8'h01, 8'h00, 8'h01, 8'h01, 8'h02, 8'h02, 8'h02,
    8'h02, 8'h01, 8'h02, 8'h02, 8'h02, 8'h00, 8'h01, 8'h02,
    8'h00, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h02,
    8'h02, 8'h01, 8'h00, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h01,
    8'h00, 8'h00, 8'h02, 8'h02, 8'h02, 8'h01, 8'h00, 8'h00,
    8'h00, 8'h00, 8'h01, 8'h00, 8'h03, 8'h02, 8'h01, 8'h01,
    8'h01, 8'h02, 8'h01, 8'h02, 8'h02, 8'h01, 8'h01, 8'h00,
    8'hFE, 8'h01, 8'h02, 8'h02, 8'h01, 8'h02, 8'h02, 8'h02,
    8'h04, 8'h02, 8'h04, 8'hFF, 8'hFB, 8'hFE, 8'h02, 8'h01,
    8'h02, 8'h01, 8'h02, 8'h02, 8'h03, 8'h01, 8'h05, 8'h06,
    8'hFF, 8'hFD, 8'h00, 8'h01, 8'h01, 8'h02, 8'h01, 8'h01,
    8'h02, 8'h02, 8'h03, 8'h07, 8'h02, 8'hFF, 8'h00, 8'h00,
    8'h02, 8'h02, 8'h02, 8'h02, 8'h01, 8'h01, 8'h04, 8'h04,
    8'h04, 8'h02, 8'h02, 8'h01, 8'hFF, 8'h02, 8'h03, 8'h02,
    8'h01, 8'h02, 8'h01, 8'h03, 8'h04, 8'h02, 8'h00, 8'h00,
    8'hFC, 8'hFF, 8'h00, 8'h01, 8'h00, 8'h02, 8'h02, 8'h03,
    8'h03, 8'h03, 8'h03, 8'h01, 8'hFD, 8'hFF, 8'h00, 8'h00,
    8'h00, 8'h02, 8'h02, 8'h01, 8'h02, 8'h03, 8'h02, 8'h01,
    8'h00, 8'hFE, 8'h00, 8'h01, 8'h01, 8'h02, 8'h01, 8'h02,
    8'h01, 8'h01, 8'h01, 8'h02, 8'h02, 8'h02, 8'h01, 8'h02,
    8'h02, 8'h01, 8'h02, 8'h01, 8'h02, 8'h00, 8'h00, 8'h00,
    8'hFD, 8'hFE, 8'hFD, 8'h02, 8'h03, 8'h02, 8'h00, 8'hFD,
    8'hFD, 8'hFF, 8'h03, 8'hFF, 8'h01, 8'hFE, 8'h00, 8'h00,
    8'h01, 8'h01, 8'h02, 8'h03, 8'h00, 8'h01, 8'hFC, 8'hFC,
    8'h04, 8'hFF, 8'hFE, 8'hFE, 8'hFF, 8'h01, 8'h00, 8'h00,
    8'h03, 8'h02, 8'h00, 8'hFE, 8'hFC, 8'h01, 8'hFF, 8'hFD,
    8'hFE, 8'hFE, 8'hFF, 8'hFF, 8'h00, 8'h01, 8'h01, 8'hFF,
    8'hFA, 8'hFC, 8'hFF, 8'h00, 8'h00, 8'hFE, 8'h00, 8'h00,
    8'hFF, 8'hFF, 8'h00, 8'h01, 8'hFE, 8'hF9, 8'hFE, 8'h02,
    8'hFE, 8'hFC, 8'hFF, 8'hFF, 8'h02, 8'h00, 8'hFF, 8'h00,
    8'h02, 8'hFD, 8'hFE, 8'hFE, 8'h00, 8'h01, 8'h00, 8'hFE,
    8'h00, 8'h02, 8'h01, 8'h00, 8'h00, 8'hFE, 8'hFD, 8'hFB,
    8'h02, 8'hFB, 8'hFE, 8'hFE, 8'hFD, 8'h01, 8'h01, 8'h00,
    8'hFC, 8'hFF, 8'hFB, 8'hFD, 8'hFE, 8'hFF, 8'hFC, 8'hFD,
    8'hFE, 8'hFD, 8'hFC, 8'h01, 8'hFF, 8'hFF, 8'hFF, 8'hFF,
    8'hFE, 8'hFF, 8'hFD, 8'hFC, 8'hFF, 8'hFF, 8'hFE, 8'hFF,
    8'h00, 8'hFF, 8'h00, 8'hFF, 8'hFD, 8'hFF, 8'h00, 8'h02,
    8'h02, 8'h01, 8'h00, 8'h00, 8'hFF, 8'hFE, 8'hFE, 8'h00,
    8'hFC, 8'hFD, 8'hFD, 8'h01, 8'hFB, 8'h00, 8'h00, 8'h00,
    8'h01, 8'hFF, 8'h01, 8'hFE, 8'h02, 8'h02, 8'hFD, 8'hFA,
    8'hFE, 8'hFF, 8'hFB, 8'hFC, 8'h01, 8'hFD, 8'hFE, 8'hFE,
    8'hFD, 8'hFC, 8'hFC, 8'hFD, 8'hFA, 8'h00, 8'h01, 8'h00,
    8'hFE, 8'hFB, 8'hFE, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFF,
    8'hFD, 8'hFC, 8'hFD, 8'h01, 8'h04, 8'h03, 8'hFF, 8'hFF,
    8'h00, 8'hFF, 8'h00, 8'h00, 8'h01, 8'h01, 8'h00, 8'h00,
    8'hFD, 8'h03, 8'hFE, 8'hFE, 8'hFE, 8'hFD, 8'hFE, 8'hFD,
    8'hFE, 8'h00, 8'h00, 8'hFF, 8'hFE, 8'hFC, 8'hFD, 8'h00,
    8'hFE, 8'hFF, 8'hFD, 8'hFE, 8'hFD, 8'hFD, 8'hFF, 8'hFF,
    8'hFB, 8'hF9, 8'hFC, 8'hFD, 8'hFF, 8'hFD, 8'hFE, 8'hFF,
    8'hFF, 8'hFE, 8'hFC, 8'hFE, 8'hFF, 8'hFC, 8'hF9, 8'hFD,
    8'hFF, 8'h00, 8'hFD, 8'hFF, 8'hFD, 8'hFD, 8'hFD, 8'hFB,
    8'hFC, 8'hFE, 8'hFB, 8'hFA, 8'h01, 8'h01, 8'hFE, 8'h00,
    8'hFE, 8'h00, 8'hFE, 8'hFB, 8'hFD, 8'hFE, 8'hFA, 8'hFE,
    8'h01, 8'h01, 8'h01, 8'hFF, 8'hFE, 8'hFE, 8'hFF, 8'hFC,
    8'hFD, 8'hFB, 8'hFF, 8'hFF, 8'h00, 8'h01, 8'hFE, 8'hFC,
    8'hFC, 8'h00, 8'hFF, 8'hFD, 8'hFD, 8'hFC, 8'h00, 8'h01,
    8'h00, 8'h01, 8'h01, 8'h00, 8'h00, 8'h02, 8'h02, 8'h00,
    8'h00, 8'h00, 8'hFC, 8'hFF, 8'h01, 8'h01, 8'hFE, 8'hFF,
    8'h01, 8'hFF, 8'h03, 8'h02, 8'h00, 8'hFD, 8'hFC, 8'hFA,
    8'hFE, 8'hFF, 8'h03, 8'hFD, 8'h00, 8'h00, 8'h02, 8'hFD,
    8'h01, 8'hFF, 8'hFF, 8'hFC, 8'hFC, 8'h03, 8'hFF, 8'hFF,
    8'h00, 8'h01, 8'hFD, 8'hFE, 8'h00, 8'h00, 8'hFC, 8'hFE,
    8'hFD, 8'hF8, 8'h02, 8'hFE, 8'hFC, 8'h01, 8'h01, 8'h00,
    8'hFF, 8'hFC, 8'hFE, 8'h01, 8'h00, 8'hFE, 8'hFA, 8'hFE,
    8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h03, 8'hFD, 8'hFD, 8'hFE,
    8'hFF, 8'hFD, 8'hF8, 8'hFA, 8'hFC, 8'hFA, 8'hFC, 8'hFE,
    8'h00, 8'h03, 8'h05, 8'h02, 8'h02, 8'h00, 8'hFD, 8'hFC,
    8'hFA, 8'hFA, 8'hFD, 8'hFB, 8'hFB, 8'hFE, 8'hFC, 8'h00,
    8'h00, 8'hFE, 8'h00, 8'hFD, 8'hFD, 8'hFC, 8'hFA, 8'hFC,
    8'hFD, 8'hFB, 8'hF9, 8'hFB, 8'hFC, 8'h02, 8'h01, 8'h00,
    8'hFD, 8'hFE, 8'hFF, 8'hFA, 8'hFA, 8'hFE, 8'hFD, 8'hFA,
    8'hFD, 8'hFC, 8'h01, 8'h00, 8'h00, 8'hFE, 8'hFE, 8'hFB,
    8'hFE, 8'hFF, 8'hFE, 8'hFC, 8'hFB, 8'h00, 8'hFF, 8'hFF,
    8'h00, 8'hFD, 8'hFC, 8'hFC, 8'hFF, 8'hFC, 8'h00, 8'h01,
    8'hFF, 8'hFB, 8'h02, 8'h00, 8'hFD, 8'h00, 8'hFC, 8'hFC,
    8'hFF, 8'hFE, 8'hF9, 8'hFD, 8'h02, 8'h01, 8'h02, 8'hFF,
    8'h00, 8'hFF, 8'hFF, 8'hFB, 8'hFC, 8'h03, 8'hFF, 8'hFD,
    8'h01, 8'h02, 8'hFF, 8'hFB, 8'hFC, 8'hFC, 8'h01, 8'h02,
    8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'h02, 8'h01, 8'h01, 8'hFF,
    8'h01, 8'h02, 8'h01, 8'h00, 8'h00, 8'hFF, 8'h00, 8'hFF,
    8'h01, 8'h04, 8'h03, 8'h02, 8'h01, 8'h02, 8'hFE, 8'h01,
    8'h00, 8'h00, 8'h01, 8'h01, 8'h01, 8'h01, 8'h02, 8'h02,
    8'hFF, 8'hFD, 8'h03, 8'hFD, 8'hFB, 8'hFD, 8'h00, 8'hFD,
    8'h00, 8'hFF, 8'hFE, 8'h00, 8'h00, 8'h00, 8'hFB, 8'hFE,
    8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'hFF,
    8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'hFF,
    8'hFF, 8'hFF, 8'hFE, 8'hFF, 8'h00, 8'hFF, 8'h00, 8'hFF,
    8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h02, 8'h01, 8'h01,
    8'hFE, 8'hFC, 8'hFC, 8'hFC, 8'hFD, 8'hFF, 8'hFF, 8'h00,
    8'hFF, 8'h02, 8'h04, 8'h02, 8'h01, 8'h00, 8'hFF, 8'hFD,
    8'hFC, 8'hFE, 8'hFE, 8'h00, 8'hFF, 8'h00, 8'h03, 8'h02,
    8'h03, 8'h01, 8'h00, 8'hFF, 8'hFF, 8'hFE, 8'hFE, 8'h00,
    8'h00, 8'hFF, 8'hFF, 8'h04, 8'h05, 8'h04, 8'h04, 8'h03,
    8'h03, 8'h01, 8'hFF, 8'h01, 8'h00, 8'hFF, 8'hFF, 8'h00,
    8'h05, 8'h06, 8'h03, 8'h01, 8'h00, 8'h02, 8'h04, 8'h02,
    8'h01, 8'h03, 8'h00, 8'hFF, 8'h00, 8'h01, 8'h04, 8'h02,
    8'h00, 8'hFE, 8'h02, 8'h02, 8'h02, 8'h01, 8'h03, 8'hFF,
    8'hFF, 8'hFF, 8'hFD, 8'hFF, 8'h01, 8'h01, 8'h02, 8'h03,
    8'h01, 8'h02, 8'h04, 8'h00, 8'h00, 8'hFF, 8'h00, 8'h00,
    8'h00, 8'hFF, 8'h02, 8'h01, 8'hFF, 8'h00, 8'h00, 8'h01,
    8'h00, 8'hFF, 8'hFF, 8'h00, 8'hFF, 8'hFE, 8'hFF, 8'h00,
    8'h00, 8'h00, 8'hFF, 8'h00, 8'h00, 8'h00, 8'hFF, 8'h00,
    8'h00, 8'h00, 8'hFF, 8'h00, 8'hFF, 8'hFE, 8'hFF, 8'h00,
    8'h00, 8'hFF, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF,
    8'h01, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF,
    8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h03, 8'h03, 8'hFE,
    8'hFE, 8'h00, 8'hFD, 8'hFF, 8'h02, 8'h01, 8'hFE, 8'hFE,
    8'h01, 8'h00, 8'hFF, 8'h01, 8'h00, 8'hFF, 8'h00, 8'hFC,
    8'hFF, 8'hFF, 8'h02, 8'h01, 8'h01, 8'h00, 8'hFF, 8'h01,
    8'h01, 8'h00, 8'h00, 8'h00, 8'hFD, 8'hFF, 8'hFD, 8'h03,
    8'hFF, 8'h02, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF,
    8'hFF, 8'hFE, 8'h00, 8'hFF, 8'h00, 8'hFF, 8'hFD, 8'hFE,
    8'hFD, 8'hFE, 8'hFD, 8'hFE, 8'hFF, 8'h00, 8'h00, 8'h01,
    8'h01, 8'hFC, 8'hFF, 8'hFE, 8'hFE, 8'hFB, 8'hFC, 8'hFD,
    8'hFD, 8'hFE, 8'h00, 8'h01, 8'h00, 8'h02, 8'h02, 8'h00,
    8'hFE, 8'hFE, 8'h00, 8'h00, 8'h01, 8'hFF, 8'hFF, 8'h00,
    8'h01, 8'h00, 8'h01, 8'h02, 8'h02, 8'h00, 8'h01, 8'h01,
    8'h03, 8'h02, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
    8'h02, 8'h03, 8'h00, 8'h02, 8'h03, 8'h03, 8'h03, 8'h02,
    8'h00, 8'hFE, 8'hFE, 8'hFF, 8'hFE, 8'h02, 8'h01, 8'h01,
    8'h00, 8'h01, 8'h02, 8'h01, 8'h00, 8'h01, 8'hFF, 8'hFE,
    8'hFF, 8'hFD, 8'hFF, 8'h04, 8'h01, 8'h01, 8'h01, 8'h00,
    8'h01, 8'h00, 8'hFF, 8'h00, 8'hFE, 8'hFC, 8'hFD, 8'hFF,
    8'h04, 8'h00, 8'h00, 8'h00, 8'hFF, 8'h02, 8'h00, 8'hFF,
    8'hFF, 8'hFD, 8'hFD, 8'hFD, 8'h00, 8'hFB, 8'hFD, 8'h00,
    8'hFE, 8'hFC, 8'hFC, 8'hFF, 8'hFD, 8'hFE, 8'hFB, 8'hFC,
    8'hFE, 8'h00, 8'hFC, 8'hFD, 8'hFF, 8'hFE, 8'h01, 8'h01,
    8'h00, 8'h00, 8'h01, 8'hFE, 8'hFC, 8'h01, 8'h00, 8'hFE,
    8'hFF, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
    8'h00, 8'h01, 8'h01, 8'hFE, 8'h01, 8'h01, 8'hFF, 8'hFE,
    8'hFE, 8'hFF, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFF,
    8'hFD, 8'h02, 8'hFE, 8'hFE, 8'hFE, 8'hFF, 8'hFF, 8'hFF,
    8'hFF, 8'hFF, 8'hFE, 8'hFD, 8'h00, 8'hFC, 8'h01, 8'hFF,
    8'h00, 8'hFF, 8'hFD, 8'hFB, 8'hFD, 8'hFE, 8'h00, 8'h00,
    8'hFF, 8'hFC, 8'h02, 8'hFE, 8'hFF, 8'hFF, 8'h01, 8'h00,
    8'h00, 8'h01, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h01, 8'h04,
    8'hFF, 8'hFF, 8'h03, 8'h04, 8'h02, 8'h02, 8'h00, 8'h01,
    8'h01, 8'h00, 8'hFF, 8'h01, 8'h03, 8'h01, 8'h01, 8'h02,
    8'h01, 8'h01, 8'h01, 8'h00, 8'h01, 8'h00, 8'h01, 8'h02,
    8'h04, 8'h02, 8'h02, 8'h01, 8'h01, 8'h01, 8'h00, 8'h00,
    8'h00, 8'h02, 8'h01, 8'h00, 8'h00, 8'h02, 8'h02, 8'h03,
    8'h00, 8'h01, 8'hFF, 8'h00, 8'h01, 8'h00, 8'h02, 8'h02,
    8'h02, 8'h02, 8'h03, 8'h05, 8'h01, 8'h00, 8'h00, 8'hFF,
    8'hFF, 8'hFE, 8'hFE, 8'h01, 8'h00, 8'h02, 8'h01, 8'h06,
    8'h03, 8'hFD, 8'hFF, 8'h00, 8'h00, 8'hFC, 8'hFE, 8'hFE,
    8'hFF, 8'h02, 8'h05, 8'h03, 8'h01, 8'hFE, 8'hFA, 8'hFD,
    8'hFE, 8'hFB, 8'hF7, 8'hF3, 8'hF6, 8'hF5, 8'hF6, 8'hFC,
    8'hFD, 8'hFE, 8'hFC, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'h02,
    8'h00, 8'h03, 8'h07, 8'hFC, 8'hFC, 8'hFB, 8'h00, 8'h00,
    8'hFC, 8'hFD, 8'h01, 8'h05, 8'h01, 8'h03, 8'h03, 8'h04,
    8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'hFE, 8'h01,
    8'h01, 8'h01, 8'h01, 8'h01, 8'h03, 8'h04, 8'h03, 8'hFE,
    8'hFA, 8'h01, 8'h00, 8'hFF, 8'h01, 8'h01, 8'h00, 8'h01,
    8'h02, 8'h01, 8'h01, 8'h01, 8'hFB, 8'hF6, 8'h00, 8'h00,
    8'h02, 8'h00, 8'h01, 8'h02, 8'h01, 8'h02, 8'h01, 8'h01,
    8'hFF, 8'hFE, 8'hFA, 8'hFB, 8'hFF, 8'h01, 8'h01, 8'h02,
    8'h01, 8'h02, 8'h00, 8'h00, 8'hFD, 8'hFD, 8'hFD, 8'hFF,
    8'h02, 8'hFF, 8'h00, 8'h00, 8'h02, 8'h01, 8'h00, 8'hFF,
    8'hFC, 8'hFD, 8'hFA, 8'hFC, 8'h00, 8'h03, 8'hFE, 8'hFD,
    8'h00, 8'hFE, 8'hFE, 8'hFD, 8'h00, 8'hFD, 8'hFD, 8'hFE,
    8'hFF, 8'h02, 8'h06, 8'h05, 8'h01, 8'h00, 8'hFD, 8'hFE,
    8'hFF, 8'hFE, 8'hFE, 8'hFF, 8'h00, 8'h02, 8'h02, 8'h05,
    8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h01, 8'h02,
    8'h03, 8'h03, 8'h05, 8'h01, 8'h02, 8'h03, 8'hFF, 8'hFE,
    8'hFF, 8'h00, 8'h01, 8'h00, 8'h02, 8'h03, 8'h04, 8'h02,
    8'h02, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h01, 8'h01, 8'h01,
    8'h01, 8'h02, 8'h04, 8'h03, 8'h02, 8'hFF, 8'hFF, 8'hFA,
    8'hFB, 8'hFE, 8'hFE, 8'h00, 8'h02, 8'h01, 8'h01, 8'h01,
    8'hFF, 8'h00, 8'hFF, 8'h04, 8'hFE, 8'hFF, 8'hFF, 8'hFF,
    8'hFF, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'hFF, 8'hFE,
    8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'hFD, 8'hFD, 8'hFD,
    8'hFE, 8'hFC, 8'hFD, 8'hFD, 8'hFF, 8'hFE, 8'hFE, 8'hFE,
    8'hFE, 8'hFE, 8'hFE, 8'hFF, 8'hFC, 8'hFA, 8'hFB, 8'hFB,
    8'hFC, 8'hFE, 8'hFF, 8'hFE, 8'hFF, 8'h02, 8'h02, 8'h01,
    8'hFF, 8'hFE, 8'hFE, 8'hFF, 8'hFE, 8'hFD, 8'hFE, 8'hFF,
    8'hFF, 8'h00, 8'h02, 8'h04, 8'h04, 8'h03, 8'h02, 8'h02,
    8'h02, 8'h00, 8'hFF, 8'hFF, 8'hFE, 8'hFE, 8'h01, 8'h04,
    8'h06, 8'h06, 8'h05, 8'h02, 8'h02, 8'h02, 8'h03, 8'h02,
    8'h00, 8'hFE, 8'hFE, 8'h00, 8'h03, 8'h03, 8'h03, 8'h00,
    8'h00, 8'h00, 8'h02, 8'h01, 8'h01, 8'hFF, 8'hFF, 8'hFE,
    8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'hFF,
    8'hFF, 8'hFE, 8'hFD, 8'hFE, 8'hFE, 8'hFF, 8'hFE, 8'h00,
    8'hFF, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hFB, 8'hFE,
    8'hFF, 8'hFE, 8'hFD, 8'hFF, 8'hFD, 8'h00, 8'h01, 8'hFE,
    8'h01, 8'h00, 8'hFE, 8'hFF, 8'hFD, 8'hFE, 8'hFE, 8'hFF,
    8'hFF, 8'hFF, 8'h00, 8'h02, 8'h02, 8'h03, 8'h01, 8'h00,
    8'hFF, 8'hFE, 8'hFF, 8'hFF, 8'hFE, 8'hFF, 8'h00, 8'h01,
    8'h02, 8'h02, 8'h03, 8'h01, 8'h00, 8'hFF, 8'hFF, 8'hFF,
    8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h00,
    8'h00, 8'hFF, 8'hFF, 8'hFE, 8'hFF, 8'h00, 8'h00, 8'h00,
    8'h01, 8'hFB, 8'hFE, 8'hFD, 8'h00, 8'hFE, 8'h01, 8'hFF,
    8'hFB, 8'h00, 8'hFD, 8'h01, 8'h03, 8'h01, 8'hFF, 8'h00,
    8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFD, 8'hFF, 8'hFA, 8'hFF,
    8'h01, 8'h00, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'h01, 8'hFF,
    8'h00, 8'h00, 8'hFF, 8'hFB, 8'h02, 8'h00, 8'hFF, 8'hFE,
    8'hFF, 8'hFF, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h03,
    8'hF7, 8'h00, 8'h01, 8'hFE, 8'hFF, 8'hFF, 8'h00, 8'h01,
    8'h02, 8'h02, 8'h02, 8'h02, 8'h01, 8'hFF, 8'hFF, 8'hFF,
    8'hFF, 8'hFE, 8'h00, 8'h02, 8'h03, 8'h02, 8'h01, 8'h01,
    8'h01, 8'hFE, 8'h02, 8'hFE, 8'hFE, 8'hFB, 8'hFD, 8'hFF,
    8'h00, 8'h02, 8'h01, 8'hFF, 8'hFE, 8'hFD, 8'hFE, 8'h01,
    8'h02, 8'h01, 8'hFC, 8'hFB, 8'hFB, 8'hFD, 8'h01, 8'h01,
    8'h00, 8'hFF, 8'h00, 8'h02, 8'hFC, 8'h00, 8'h00, 8'hFD,
    8'hFC, 8'hFB, 8'hFD, 8'hFE, 8'hFF, 8'h01, 8'h01, 8'h02,
    8'h01, 8'hFA, 8'hFF, 8'h01, 8'h00, 8'h00, 8'hFF, 8'hFE,
    8'hFF, 8'h01, 8'h01, 8'h01, 8'h02, 8'h02, 8'hFB, 8'hFE,
    8'h01, 8'h00, 8'hFF, 8'h00, 8'h00, 8'h02, 8'h01, 8'h02,
    8'h02, 8'h01, 8'h02, 8'hFE, 8'hFF, 8'h02, 8'h01, 8'h00,
    8'h03, 8'h01, 8'h02, 8'h02, 8'h03, 8'h00, 8'h00, 8'h01,
    8'hFF, 8'h00, 8'hFD, 8'h01, 8'h02, 8'h02, 8'h04, 8'h02,
    8'h02, 8'h03, 8'h02, 8'hFC, 8'hF9, 8'hFE, 8'hFE, 8'h00,
    8'h02, 8'h03, 8'h00, 8'hFE, 8'hFE, 8'h01, 8'h01, 8'h02,
    8'h02, 8'hFA, 8'hFB, 8'hFF, 8'h02, 8'h00, 8'h00, 8'hFF,
    8'h01, 8'h01, 8'h01, 8'h00, 8'h00, 8'h01, 8'h02, 8'hFE,
    8'h01, 8'h00, 8'hFF, 8'h00, 8'h01, 8'h02, 8'h01, 8'hFF,
    8'hFE, 8'hFF, 8'hFF, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00,
    8'h01, 8'hFF, 8'hFF, 8'h00, 8'hFF, 8'h00, 8'hFE, 8'hFF,
    8'hFF, 8'hF7, 8'h01, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF,
    8'hFF, 8'h01, 8'h01, 8'hFF, 8'hFE, 8'hF9, 8'hF9, 8'h01,
    8'hFD, 8'hFF, 8'h00, 8'hFF, 8'h02, 8'h01, 8'h01, 8'h02,
    8'h02, 8'h00, 8'hFD, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF,
    8'hFF, 8'h00, 8'hFF, 8'h00, 8'h00, 8'h01, 8'h02, 8'h02,
    8'h01, 8'h01, 8'h00, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFD,
    8'hFF, 8'h00, 8'h00, 8'hFF, 8'h01, 8'h01, 8'h03, 8'h01,
    8'h00, 8'hFF, 8'hFE, 8'hFF, 8'h00, 8'h01, 8'h00, 8'hFE,
    8'hFE, 8'hFE, 8'hFD, 8'h02, 8'h01, 8'h00, 8'hFF, 8'hFF,
    8'hFF, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFE, 8'hFB,
    8'h02, 8'h01, 8'h02, 8'h01, 8'hFF, 8'hFF, 8'hFF, 8'hFF,
    8'h00, 8'hFF, 8'h00, 8'hF8, 8'hFF, 8'h04, 8'h00, 8'h02,
    8'h03, 8'h03, 8'h01, 8'h02, 8'h02, 8'h01, 8'h00, 8'hFF,
    8'hFA, 8'hFC, 8'h04, 8'h01, 8'h03, 8'h01, 8'hFF, 8'hFE,
    8'h00, 8'h02, 8'h03, 8'hFE, 8'hF9, 8'hFC, 8'hFD, 8'h00,
    8'hFF, 8'hFC, 8'hFC, 8'hFD, 8'hFF, 8'hFC, 8'hFC, 8'hFD,
    8'hFE, 8'hFF, 8'h00, 8'h00, 8'h03, 8'h04, 8'h02, 8'h01,
    8'h02, 8'h04, 8'h06, 8'h02, 8'h02, 8'h00, 8'hFC, 8'hFD,
    8'hFD, 8'h01, 8'h02, 8'h01, 8'h02, 8'h04, 8'h05, 8'h02,
    8'h01, 8'h02, 8'h02, 8'h01, 8'hFB, 8'hF7, 8'h02, 8'h01,
    8'h02, 8'h02, 8'h03, 8'h02, 8'h01, 8'h00, 8'hFE, 8'hFE,
    8'hFC, 8'hFD, 8'hFD, 8'h00, 8'h00, 8'h02, 8'h01, 8'h02,
    8'h01, 8'hFF, 8'h00, 8'hFE, 8'hFD, 8'hFE, 8'hFC, 8'hF7,
    8'h03, 8'h00, 8'h00, 8'h00, 8'hFF, 8'h00, 8'h01, 8'h00,
    8'h00, 8'hFF, 8'h00, 8'h01, 8'hFB, 8'hFF, 8'h00, 8'hFF,
    8'h01, 8'h00, 8'h01, 8'h03, 8'h01, 8'h02, 8'h02, 8'hFF,
    8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'h03, 8'h02, 8'h02,
    8'h04, 8'h03, 8'h03, 8'h00, 8'hFE, 8'hFB, 8'hFB, 8'h02,
    8'h00, 8'h03, 8'h02, 8'h03, 8'h05, 8'h05, 8'h03, 8'h01,
    8'hFF, 8'hFD, 8'hFB, 8'hFD, 8'h01, 8'h03, 8'h04, 8'h02,
    8'h02, 8'h04, 8'h02, 8'h03, 8'h00, 8'hFE, 8'hFD, 8'hFC,
    8'hFA, 8'h01, 8'h02, 8'h03, 8'h03, 8'h01, 8'h00, 8'h01,
    8'h00, 8'hFD, 8'hFE, 8'hFC, 8'hFE, 8'hFF, 8'h04, 8'h00,
    8'h02, 8'h01, 8'h02, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFE,
    8'h00, 8'h02, 8'h00, 8'h03, 8'h02, 8'h02, 8'h01, 8'h01,
    8'h02, 8'h00, 8'h00, 8'h01, 8'hFE, 8'h00, 8'h01, 8'hFC,
    8'h01, 8'h01, 8'h01, 8'h02, 8'h01, 8'h02, 8'h01, 8'h01,
    8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h00,
    8'h01, 8'h01, 8'h01, 8'h00, 8'h00, 8'h01, 8'h00, 8'hFF,
    8'h00, 8'h01, 8'h01, 8'h01, 8'h00, 8'hFF, 8'h00, 8'h00,
    8'hFE, 8'h00, 8'hFE, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01,
    8'h01, 8'h00, 8'hFF, 8'hFE, 8'h00, 8'hFE, 8'hFF, 8'hFF,
    8'h01, 8'h02, 8'h01, 8'h00, 8'h01, 8'h00, 8'h00, 8'hFD,
    8'hFE, 8'h00, 8'h02, 8'h01, 8'hFE, 8'h00, 8'h01, 8'h01,
    8'h01, 8'h00, 8'h01, 8'hFF, 8'hFB, 8'hFF, 8'hFF, 8'h02,
    8'hFF, 8'hFB, 8'hFE, 8'h00, 8'h01, 8'h01, 8'h01, 8'hFE,
    8'hFC, 8'hFC, 8'hFE, 8'hFF, 8'hFF, 8'hF8, 8'hFD, 8'hFF,
    8'h01, 8'h01, 8'h01, 8'h01, 8'h00, 8'hFF, 8'hFF, 8'hFF,
    8'hFF, 8'h02, 8'h00, 8'h01, 8'h00, 8'h02, 8'h00, 8'h01,
    8'h01, 8'h01, 8'h02, 8'h01, 8'h00, 8'hFF, 8'h00, 8'hFE,
    8'h00, 8'h01, 8'h00, 8'h02, 8'h02, 8'h00, 8'h01, 8'h02,
    8'h02, 8'h03, 8'h01, 8'hFF, 8'hFE, 8'hFE, 8'h00, 8'h01,
    8'h02, 8'h01, 8'h01, 8'h01, 8'h02, 8'h03, 8'h03, 8'h02,
    8'h01, 8'hFE, 8'hFE, 8'hFF, 8'h00, 8'h01, 8'h01, 8'h01,
    8'h01, 8'h01, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00,
    8'h00, 8'h02, 8'h01, 8'h00, 8'h01, 8'h01, 8'h01, 8'h01,
    8'h03, 8'h01, 8'h02, 8'h01, 8'h01, 8'h02, 8'h00, 8'h01,
    8'h01, 8'h00, 8'h00, 8'hFB, 8'hFB, 8'hF8, 8'hF9, 8'hFD,
    8'hFB, 8'hFA, 8'hF6, 8'hFD, 8'hFC, 8'hFD, 8'hFF, 8'h01,
    8'hFE, 8'hFD, 8'hFE, 8'hFF, 8'h01, 8'h02, 8'h00, 8'h03,
    8'h02, 8'h02, 8'hFF, 8'hFE, 8'hFB, 8'h00, 8'h01, 8'hFE,
    8'hFF, 8'h01, 8'h02, 8'h02, 8'h01, 8'h03, 8'h03, 8'hFF,
    8'hFE, 8'hFF, 8'hFE, 8'h01, 8'h00, 8'hFF, 8'hFF, 8'h01,
    8'h02, 8'h02, 8'h03, 8'h01, 8'h03, 8'h00, 8'hFF, 8'h00,
    8'h00, 8'h01, 8'h01, 8'hFE, 8'h01, 8'h03, 8'h01, 8'h01,
    8'hFF, 8'hFE, 8'h00, 8'hFD, 8'h01, 8'h02, 8'h02, 8'h01,
    8'hFC, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFD, 8'hFE, 8'hFD,
    8'h01, 8'h01, 8'h02, 8'h02, 8'h00, 8'hFD, 8'hFF, 8'h00,
    8'h01, 8'hFF, 8'hFD, 8'hFF, 8'hFF, 8'h02, 8'hFF, 8'h01,
    8'h00, 8'hFF, 8'hFF, 8'h01, 8'h01, 8'h01, 8'hFF, 8'hFC,
    8'hFE, 8'hFF, 8'h01, 8'h00, 8'h00, 8'hFF, 8'h00, 8'hFF,
    8'h01, 8'h01, 8'h00, 8'h00, 8'hFE, 8'hFD, 8'h01, 8'hFF,
    8'h00, 8'h01, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFE,
    8'hFF, 8'hFC, 8'hFC, 8'hFE, 8'hFE, 8'hFE, 8'h01, 8'h00,
    8'h00, 8'h00, 8'h00, 8'hFE, 8'hFE, 8'hFF, 8'hFF, 8'hFC,
    8'hFE, 8'hF6, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFE,
    8'hFE, 8'h01, 8'h02, 8'hFF, 8'hFE, 8'hFF, 8'h02, 8'h00,
    8'hFD, 8'hFD, 8'hFB, 8'hFD, 8'hFE, 8'hFF, 8'hFE, 8'hFF,
    8'hFC, 8'hFF, 8'hFF, 8'hFD, 8'hFB, 8'hFC, 8'hFB, 8'hFB,
    8'hFD, 8'h00, 8'hFF, 8'h00, 8'h01, 8'hFD, 8'hFD, 8'hFE,
    8'hFD, 8'hFE, 8'h00, 8'h00, 8'h01, 8'h01, 8'h01, 8'h01,
    8'h01, 8'h01, 8'h01, 8'hFF, 8'hFE, 8'h00, 8'h02, 8'h02,
    8'h01, 8'hFF, 8'hFE, 8'h00, 8'h00, 8'hFF, 8'h00, 8'h01,
    8'h03, 8'hFF, 8'h01, 8'h01, 8'h00, 8'hFF, 8'hFE, 8'hFE,
    8'hFF, 8'h00, 8'h01, 8'h01, 8'hFE, 8'h00, 8'hFF, 8'hFF,
    8'hFF, 8'h00, 8'h01, 8'hFF, 8'h00, 8'h01, 8'h00, 8'h01,
    8'h00, 8'hFD, 8'hFA, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h02,
    8'h02, 8'h03, 8'h01, 8'h00, 8'h01, 8'h01, 8'hFF, 8'hFC,
    8'hFF, 8'h02, 8'hFE, 8'h00, 8'h01, 8'h01, 8'h02, 8'h00,
    8'h01, 8'h02, 8'hFF, 8'h00, 8'hFD, 8'h00, 8'hFE, 8'hFD,
    8'h00, 8'h01, 8'h01, 8'h02, 8'h02, 8'h00, 8'h01, 8'h00,
    8'hFD, 8'hFF, 8'hFE, 8'hFF, 8'h01, 8'hFE, 8'hFF, 8'h00,
    8'h01, 8'h01, 8'h00, 8'hFF, 8'h00, 8'hFF, 8'hFF, 8'hFE,
    8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD,
    8'hFC, 8'hFB, 8'h00, 8'hFC, 8'hFE, 8'hFD, 8'h01, 8'h00,
    8'h00, 8'hFF, 8'hFF, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'hFF,
    8'hFF, 8'hFE, 8'hFD, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'h02,
    8'h02, 8'h01, 8'h00, 8'h00, 8'h03, 8'h00, 8'hFF, 8'h01,
    8'hFE, 8'h00, 8'hFE, 8'hFF, 8'h01, 8'h03, 8'hFD, 8'hFE,
    8'hFC, 8'hFC, 8'h00, 8'h00, 8'hFE, 8'hFB, 8'hFD, 8'hFC,
    8'hFD, 8'hFC, 8'hF8, 8'hF8, 8'hFB, 8'hFC, 8'hFD, 8'h00,
    8'hFD, 8'hFC, 8'hFB, 8'hFA, 8'hFC, 8'hFA, 8'hFC, 8'hFA,
    8'hFC, 8'hFD, 8'hFB, 8'hFD, 8'hFE, 8'hFD, 8'hFC, 8'hFF,
    8'h01, 8'hFE, 8'hFF, 8'hFD, 8'hFB, 8'hFD, 8'hFC, 8'h01,
    8'h02, 8'hFE, 8'hFF, 8'h01, 8'hFF, 8'hFE, 8'hFF, 8'hFB,
    8'hF9, 8'hF7, 8'hF6, 8'hFA, 8'hFD, 8'hFF, 8'hFF, 8'hFD,
    8'h00, 8'hFF, 8'hFD, 8'hFB, 8'hFB, 8'hFA, 8'hFA, 8'hF9,
    8'hFB, 8'hFD, 8'hFF, 8'h02, 8'h00, 8'hFF, 8'hFC, 8'hFF,
    8'hFF, 8'hFD, 8'hF9, 8'hFD, 8'hFD, 8'hFD, 8'hFD, 8'hFD,
    8'hFC, 8'hFD, 8'hFE, 8'h00, 8'hFF, 8'h00, 8'h02, 8'hFF,
    8'hFC, 8'h00, 8'h02, 8'h01, 8'h02, 8'hFE, 8'h01, 8'h02,
    8'h01, 8'h01, 8'h01, 8'h03, 8'h01, 8'h00, 8'h00, 8'h00,
    8'h00, 8'h00, 8'hFE, 8'hFD, 8'h00, 8'h00, 8'h00, 8'h00,
    8'h01, 8'h01, 8'h02, 8'h01, 8'h02, 8'h02, 8'h01, 8'hFD,
    8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFE, 8'hFF, 8'h00, 8'hFF,
    8'h02, 8'h02, 8'hFF, 8'hFF, 8'hFC, 8'hFF, 8'hFE, 8'hFD,
    8'hFD, 8'hFC, 8'hFB, 8'hFE, 8'h01, 8'h02, 8'h05, 8'h02,
    8'hFE, 8'hFC, 8'hFD, 8'hF9, 8'hFD, 8'hFD, 8'hFC, 8'hFD,
    8'hFE, 8'hFF, 8'h01, 8'h01, 8'h01, 8'hFF, 8'hFD, 8'hFE,
    8'h02, 8'hFF, 8'hFE, 8'h00, 8'hFF, 8'h01, 8'h00, 8'h00,
    8'h00, 8'h00, 8'h01, 8'hFC, 8'h00, 8'h00, 8'h00, 8'h00,
    8'h00, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00,
    8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01,
    8'h00, 8'h00, 8'h00, 8'h01, 8'hFF, 8'hFF, 8'h00, 8'h00,
    8'hFF, 8'hFE, 8'hFF, 8'h01, 8'h05, 8'h04, 8'h05, 8'h06,
    8'h06, 8'h01, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFC, 8'hFC,
    8'hFE, 8'h02, 8'h04, 8'h05, 8'h06, 8'h05, 8'h01, 8'h00,
    8'h00, 8'h00, 8'hFE, 8'hFC, 8'hFA, 8'hFD, 8'hFE, 8'hFF,
    8'h02, 8'h03, 8'h03, 8'h02, 8'h00, 8'h00, 8'h00, 8'hFF,
    8'hFD, 8'hFE, 8'hFD, 8'hFE, 8'h00, 8'h00, 8'hFE, 8'h01,
    8'h01, 8'h01, 8'h00, 8'h00, 8'h00, 8'h01, 8'hFF, 8'hFE,
    8'h00, 8'h01, 8'hFD, 8'hFC, 8'hFE, 8'h00, 8'h00, 8'hFF,
    8'h00, 8'h01, 8'h02, 8'hFF, 8'h00, 8'h02, 8'h01, 8'hFC,
    8'hFB, 8'hFC, 8'hFD, 8'h00, 8'h00, 8'hFF, 8'h00, 8'h01,
    8'h02, 8'h01, 8'h00, 8'h00, 8'hFF, 8'hFD, 8'hFD, 8'hFE,
    8'h00, 8'h00, 8'h00, 8'h01, 8'h01, 8'h02, 8'h01, 8'h01,
    8'h01, 8'h00, 8'h00, 8'hFE, 8'hFF, 8'hFE, 8'hFF, 8'hFF,
    8'h02, 8'h01, 8'h01, 8'h00, 8'h02, 8'h01, 8'h01, 8'h01,
    8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF,
    8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h00, 8'h00, 8'h01,
    8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'hFF,
    8'h00, 8'h00, 8'h00, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'h00,
    8'hFE, 8'hFF, 8'hFC, 8'hFD, 8'hFF, 8'h01, 8'h01, 8'h00,
    8'hFD, 8'hFE, 8'hFE, 8'hFD, 8'hFD, 8'hFE, 8'h00, 8'h00,
    8'h00, 8'h01, 8'h03, 8'h01, 8'h01, 8'h01, 8'h02, 8'h01,
    8'hFE, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'h00, 8'h01,
    8'h00, 8'h01, 8'h03, 8'h03, 8'hFD, 8'hFE, 8'h00, 8'h01,
    8'h00, 8'h00, 8'hFE, 8'hFD, 8'hFE, 8'h00, 8'h00, 8'h02,
    8'h03, 8'hFB, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFD,
    8'hFC, 8'hFC, 8'hFB, 8'hFC, 8'h01, 8'h04, 8'hFC, 8'h01,
    8'hFE, 8'hFF, 8'h00, 8'h01, 8'hFF, 8'hFD, 8'hFC, 8'hFA,
    8'hF9, 8'hFD, 8'h00, 8'hFF, 8'hFE, 8'hFD, 8'hFD, 8'h00,
    8'h01, 8'h01, 8'hFE, 8'hFF, 8'hFD, 8'hFC, 8'hFB, 8'hFE,
    8'hFA, 8'hFE, 8'hFD, 8'hFB, 8'hFF, 8'h00, 8'hFF, 8'hFF,
    8'hFF, 8'hFF, 8'hFF, 8'h00, 8'hFC, 8'hFB, 8'h00, 8'h01,
    8'hFD, 8'hFE, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00,
    8'h01, 8'hFE, 8'h01, 8'h00, 8'h01, 8'hFF, 8'h00, 8'h00,
    8'hFF, 8'h00, 8'h00, 8'h01, 8'h00, 8'h02, 8'h03, 8'h00,
    8'h00, 8'h00, 8'h01, 8'h00, 8'h01, 8'h01, 8'h00, 8'h01,
    8'h02, 8'h02, 8'h03, 8'h04, 8'hFD, 8'h01, 8'hFF, 8'h01,
    8'h01, 8'h01, 8'h01, 8'h02, 8'h01, 8'h01, 8'h00, 8'h02,
    8'h02, 8'h01, 8'hFE, 8'hFE, 8'hFF, 8'hFE, 8'h00, 8'h02,
    8'h02, 8'h02, 8'h02, 8'h01, 8'h05, 8'hFD, 8'hFB, 8'h00,
    8'h00, 8'hFD, 8'h00, 8'h00, 8'hFF, 8'h01, 8'h00, 8'h01,
    8'h01, 8'hFF, 8'hFE, 8'hFC, 8'hFF, 8'h00, 8'hFF, 8'h02,
    8'h00, 8'hFF, 8'hFF, 8'h00, 8'hFF, 8'hFE, 8'hFF, 8'h01,
    8'hFE, 8'h01, 8'h00, 8'h00, 8'h01, 8'h00, 8'hFF, 8'hFF,
    8'h01, 8'h00, 8'h02, 8'h01, 8'h00, 8'hF9, 8'h01, 8'hFF,
    8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFE, 8'hFE, 8'h01, 8'h02,
    8'h03, 8'h04, 8'hF8, 8'h00, 8'h00, 8'hFE, 8'hFF, 8'hFF,
    8'hFF, 8'hFE, 8'hFC, 8'hFF, 8'hFF, 8'h02, 8'h04, 8'hFC,
    8'hFE, 8'hFD, 8'hFD, 8'hFF, 8'hFF, 8'h00, 8'hFF, 8'hFE,
    8'hFE, 8'hFF, 8'h00, 8'h03, 8'h00, 8'hFE, 8'hFF, 8'hFD,
    8'hFE, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'h00, 8'h00,
    8'h05, 8'hFE, 8'hFD, 8'h01, 8'hFF, 8'h00, 8'hFF, 8'hFF,
    8'h00, 8'hFF, 8'hFE, 8'hFF, 8'h01, 8'h00, 8'hFF, 8'h02,
    8'h01, 8'h00, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFE,
    8'h00, 8'hFE, 8'h01, 8'hFE, 8'h01, 8'hFF, 8'hFF, 8'hFF,
    8'hFF, 8'h01, 8'h01, 8'h00, 8'h00, 8'hFF, 8'hFC, 8'hFF,
    8'hFD, 8'h01, 8'hFF, 8'h01, 8'hFF, 8'hFF, 8'h00, 8'h00,
    8'h01, 8'h00, 8'h01, 8'hFD, 8'hFF, 8'h01, 8'hFF, 8'h02,
    8'h01, 8'h01, 8'h01, 8'h02, 8'h01, 8'h02, 8'hFF, 8'h05,
    8'hFD, 8'h01, 8'hFF, 8'hFD, 8'hFD, 8'hFE, 8'hFB, 8'h00,
    8'hFF, 8'h01, 8'hFF, 8'h00, 8'h03, 8'hFA, 8'hFB, 8'h00,
    8'h00, 8'hFE, 8'hFD, 8'hFE, 8'hFF, 8'hFC, 8'hFF, 8'hFF,
    8'hFF, 8'h00, 8'hFF, 8'h00, 8'hFA, 8'h00, 8'hFB, 8'hFD,
    8'hFC, 8'hFB, 8'hFE, 8'hFE, 8'h00, 8'hFF, 8'hFF, 8'h01,
    8'hFF, 8'h01, 8'h00, 8'hFD, 8'hFC, 8'hFF, 8'hFE, 8'hFE,
    8'hFF, 8'hFE, 8'hFE, 8'h00, 8'h03, 8'hFF, 8'hFD, 8'hFE,
    8'hFD, 8'hFE, 8'hFE, 8'h01, 8'h00, 8'h01, 8'h01, 8'h02,
    8'h00, 8'h01, 8'h03, 8'hF9, 8'hFF, 8'hFD, 8'h01, 8'h01,
    8'h01, 8'h02, 8'h03, 8'h05, 8'h03, 8'h02, 8'h04, 8'h02,
    8'hFA, 8'h00, 8'h01, 8'h00, 8'h00, 8'h01, 8'h03, 8'h04,
    8'h05, 8'h04, 8'h04, 8'h06, 8'h07, 8'h01, 8'h00, 8'h03,
    8'h03, 8'h02, 8'h03, 8'h02, 8'h03, 8'h03, 8'h03, 8'h03,
    8'hFF, 8'h04, 8'hFF, 8'h02, 8'h03, 8'h05, 8'h03, 8'h03,
    8'h02, 8'h00, 8'h01, 8'h02, 8'h02, 8'hFF, 8'hFE, 8'hFF,
    8'h02, 8'h01, 8'h03, 8'h04, 8'h01, 8'h01, 8'h01, 8'h01,
    8'h01, 8'h00, 8'hFE, 8'hFE, 8'h00, 8'h02, 8'h03, 8'h02,
    8'h00, 8'hFF, 8'h01, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFF,
    8'hFC, 8'hFD, 8'h01, 8'h01, 8'h03, 8'h01, 8'h00, 8'h01,
    8'h00, 8'hFF, 8'hFE, 8'h00, 8'h00, 8'hFF, 8'h01, 8'h01,
    8'h00, 8'h03, 8'h02, 8'h01, 8'h00, 8'hFF, 8'hFF, 8'hFF,
    8'hFF, 8'h02, 8'h03, 8'h00, 8'hFD, 8'hFF, 8'h02, 8'h02,
    8'h02, 8'h01, 8'h01, 8'h00, 8'hFF, 8'h01, 8'h01, 8'hFF,
    8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF,
    8'h00, 8'hFF, 8'hFF, 8'h01, 8'h01, 8'h00, 8'h00, 8'h00,
    8'hFF, 8'hFE, 8'h00, 8'h01, 8'h04, 8'h02, 8'h00, 8'h01,
    8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'h01, 8'hFE,
    8'h02, 8'h04, 8'h05, 8'h02, 8'h00, 8'hFF, 8'h00, 8'h00,
    8'h00, 8'h00, 8'h00, 8'h02, 8'h03, 8'h04, 8'h05, 8'h06,
    8'h04, 8'h02, 8'h03, 8'h00, 8'h00, 8'h00, 8'hFF, 8'h00,
    8'hFF, 8'h04, 8'h03, 8'h07, 8'h05, 8'h05, 8'h04, 8'h00,
    8'hFF, 8'h00, 8'h00, 8'hFE, 8'h00, 8'hFE, 8'hFE, 8'h01,
    8'h04, 8'h03, 8'h00, 8'hFE, 8'hFD, 8'h00, 8'h01, 8'h01,
    8'hFD, 8'hFE, 8'hFC, 8'hFA, 8'h02, 8'h02, 8'hFF, 8'hFC,
    8'hFE, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFE, 8'hFD, 8'hF9,
    8'hFD, 8'h00, 8'hFD, 8'hFE, 8'h01, 8'h01, 8'h00, 8'h00,
    8'h00, 8'h01, 8'h00, 8'hFA, 8'hF9, 8'hFA, 8'hFD, 8'hFF,
    8'h00, 8'h02, 8'h01, 8'h01, 8'h00, 8'hFF, 8'h00, 8'hFF,
    8'hFE, 8'hFA, 8'hF9, 8'hFD, 8'h02, 8'h02, 8'h01, 8'h01,
    8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFD, 8'hFB,
    8'hFF, 8'h01, 8'h01, 8'h01, 8'hFF, 8'h00, 8'h00, 8'h00,
    8'h00, 8'h00, 8'h01, 8'h02, 8'hFF, 8'hFF, 8'h00, 8'h00,
    8'h00, 8'h00, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00,
    8'h00, 8'h00, 8'h00, 8'h01, 8'h01, 8'h00, 8'h00, 8'h00,
    8'h00, 8'h00, 8'h00, 8'h05, 8'h05, 8'h06, 8'h04, 8'h03,
    8'h05, 8'h02, 8'h04, 8'h04, 8'h03, 8'h00, 8'hFE, 8'h01,
    8'h02, 8'h02, 8'h03, 8'h02, 8'h01, 8'hFF, 8'h00, 8'h02,
    8'h02, 8'h01, 8'hFE, 8'hFE, 8'h02, 8'h01, 8'h03, 8'h01,
    8'h00, 8'h00, 8'h00, 8'hFF, 8'h00, 8'hFF, 8'h00, 8'h00,
    8'hFD, 8'h03, 8'h00, 8'h01, 8'h01, 8'hFF, 8'hFF, 8'hFE,
    8'hFD, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'hFD, 8'h02, 8'h00,
    8'h02, 8'h01, 8'hFF, 8'hFF, 8'hFD, 8'hFC, 8'hFD, 8'hFD,
    8'hFC, 8'hFB, 8'hFC, 8'hFF, 8'h02, 8'h01, 8'h01, 8'h01,
    8'h00, 8'hFF, 8'hFD, 8'hFE, 8'hFF, 8'h00, 8'hFD, 8'hFD,
    8'hFE, 8'h02, 8'h01, 8'h01, 8'h02, 8'h01, 8'h01, 8'hFE,
    8'hFF, 8'h00, 8'h02, 8'hFF, 8'hFC, 8'hFC, 8'h01, 8'h01,
    8'h02, 8'h02, 8'h02, 8'h03, 8'h00, 8'h00, 8'h01, 8'h02,
    8'h03, 8'hFD, 8'hFF, 8'hFF, 8'h01, 8'h01, 8'h01, 8'h01,
    8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'hFB, 8'hFD,
    8'hFE, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00,
    8'hFF, 8'hFF, 8'h01, 8'hFE, 8'hFE, 8'hFF, 8'hFF, 8'h00,
    8'h00, 8'hFF, 8'h01, 8'h00, 8'h00, 8'h00, 8'hFD, 8'hFF,
    8'h00, 8'hFB, 8'hF8, 8'hFE, 8'hFF, 8'hFF, 8'hFE, 8'h01,
    8'h01, 8'h03, 8'hFD, 8'hFC, 8'hFD, 8'hFF, 8'hFF, 8'hFD,
    8'hFB, 8'hF8, 8'h00, 8'hFD, 8'h00, 8'hFE, 8'hFB, 8'hFC,
    8'hFF, 8'h00, 8'h01, 8'hFF, 8'h03, 8'h04, 8'h02, 8'h02,
    8'h03, 8'h01, 8'hFF, 8'h02, 8'h01, 8'h02, 8'h02, 8'hFE,
    8'h01, 8'h01, 8'h03, 8'h02, 8'hFF, 8'hFF, 8'h00, 8'h00,
    8'h00, 8'h00, 8'h01, 8'h03, 8'hFC, 8'h02, 8'h01, 8'h01,
    8'hFE, 8'hFD, 8'hFE, 8'hFE, 8'hFE, 8'hFF, 8'hFE, 8'hFD,
    8'h02, 8'hFD, 8'h01, 8'h01, 8'hFF, 8'h00, 8'hFF, 8'hFF,
    8'hFF, 8'hFD, 8'hFE, 8'h00, 8'hFE, 8'hFA, 8'hFC, 8'hFE,
    8'h00, 8'h01, 8'h01, 8'h01, 8'h02, 8'h02, 8'h00, 8'h00,
    8'h01, 8'h02, 8'h00, 8'hFB, 8'h00, 8'h00, 8'h02, 8'hFF,
    8'h01, 8'h00, 8'h02, 8'h02, 8'h01, 8'h01, 8'h01, 8'h01,
    8'hFB, 8'h01, 8'h00, 8'h01, 8'hFE, 8'hFF, 8'h02, 8'h04,
    8'h02, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFC, 8'h02, 8'h01,
    8'h01, 8'h00, 8'hFD, 8'h02, 8'h03, 8'h02, 8'h01, 8'h00,
    8'hFE, 8'hFE, 8'hFD, 8'h02, 8'hFF, 8'hFF, 8'h00, 8'hFF,
    8'hFF, 8'h01, 8'h00, 8'h01, 8'h01, 8'h02, 8'hFD, 8'hFF,
    8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01,
    8'h02, 8'h01, 8'h03, 8'hFB, 8'hFF, 8'hFD, 8'hFD, 8'hFE,
    8'hFD, 8'hFE, 8'h02, 8'h02, 8'h03, 8'h03, 8'h00, 8'hFB,
    8'h00, 8'h00, 8'hFB, 8'h00, 8'h02, 8'hFC, 8'hFA, 8'hFB,
    8'hFA, 8'hFF, 8'hFA, 8'hFB, 8'hFE, 8'h01, 8'h02, 8'h00,
    8'hFE, 8'hFC, 8'hFF, 8'hFC, 8'hFB, 8'hFD, 8'hFA, 8'hFE,
    8'h00, 8'h01, 8'h01, 8'h01, 8'h02, 8'h04, 8'h04, 8'h01,
    8'h00, 8'hFD, 8'hFD, 8'h04, 8'h05, 8'h04, 8'h01, 8'h00,
    8'h00, 8'h00, 8'h04, 8'h00, 8'hFC, 8'hFA, 8'hFC, 8'hFD,
    8'hFE, 8'hFF, 8'h02, 8'hFF, 8'hFD, 8'hFB, 8'h00, 8'hFE,
    8'hFD, 8'hFA, 8'hFA, 8'hFB, 8'hFD, 8'hFF, 8'hFF, 8'hFF,
    8'h01, 8'hFF, 8'hFC, 8'hFE, 8'hFF, 8'hFE, 8'hF8, 8'hFA,
    8'hFC, 8'hFD, 8'hFF, 8'h01, 8'h02, 8'h03, 8'h00, 8'hFC,
    8'hFE, 8'hFE, 8'hFC, 8'hF7, 8'hF9, 8'hFA, 8'hFD, 8'hFF,
    8'h03, 8'h03, 8'hFF, 8'hF9, 8'hFB, 8'hFC, 8'hFD, 8'hFD,
    8'hF8, 8'hFB, 8'hFC, 8'hFF, 8'h02, 8'h03, 8'h02, 8'hFE,
    8'hFA, 8'hFB, 8'hFF, 8'hFD, 8'hFB, 8'hFA, 8'hFB, 8'hFE,
    8'h03, 8'h02, 8'h02, 8'h01, 8'h01, 8'hF9, 8'hFB, 8'hFF,
    8'h00, 8'hFD, 8'hFC, 8'hFD, 8'h00, 8'h02, 8'h01, 8'h01,
    8'h00, 8'h00, 8'hFA, 8'hFB, 8'h00, 8'hFF, 8'hFF, 8'hFF,
    8'hFF, 8'hFE, 8'h00, 8'h01, 8'h01, 8'hFE, 8'h00, 8'hFE,
    8'hFE, 8'hFE, 8'hFF, 8'h00, 8'h00, 8'h02, 8'h01, 8'h01,
    8'h01, 8'hFF, 8'hFD, 8'h00, 8'h01, 8'hFC, 8'hFD, 8'h01,
    8'hFF, 8'h01, 8'h02, 8'h02, 8'h02, 8'h01, 8'hFE, 8'hFD,
    8'hFF, 8'h02, 8'hFF, 8'hF8, 8'hFB, 8'h00, 8'h00, 8'h01,
    8'h00, 8'h00, 8'hFF, 8'h01, 8'hFE, 8'hF9, 8'hFC, 8'hFF,
    8'hFF, 8'hFC, 8'hFA, 8'hF8, 8'hFF, 8'h00, 8'h00, 8'h00,
    8'hFD, 8'hFA, 8'hFC, 8'hFF, 8'h00, 8'h01, 8'h00, 8'h00,
    8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00,
    8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h02, 8'h01,
    8'h01, 8'h01, 8'h01, 8'h00, 8'h00, 8'h01, 8'h00, 8'h01,
    8'h00, 8'h01, 8'hFF, 8'hFE, 8'h00, 8'h01, 8'h00, 8'h01,
    8'h00, 8'h01, 8'h01, 8'h01, 8'h00, 8'hFE, 8'hFD, 8'hFE,
    8'hFE, 8'h00, 8'hFF, 8'hFE, 8'hFF, 8'h00, 8'h01, 8'h00,
    8'h00, 8'h00, 8'hFE, 8'hFE, 8'hFF, 8'h00, 8'h00, 8'hFD,
    8'hFE, 8'hFF, 8'hFF, 8'h01, 8'h01, 8'h00, 8'h00, 8'h00,
    8'h00, 8'h02, 8'h02, 8'h01, 8'h00, 8'h00, 8'h01, 8'h01,
    8'h00, 8'h00, 8'h00, 8'h02, 8'h01, 8'h03, 8'h06, 8'h06,
    8'h02, 8'h02, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'h00, 8'h00,
    8'h02, 8'h04, 8'h05, 8'h08, 8'h04, 8'hFF, 8'h01, 8'h02,
    8'h03, 8'h00, 8'h02, 8'h00, 8'h01, 8'h01, 8'h02, 8'h04,
    8'h05, 8'h00, 8'hFF, 8'hFF, 8'h02, 8'h02, 8'h02, 8'h01,
    8'h00, 8'h00, 8'h02, 8'h02, 8'h02, 8'h02, 8'h01, 8'hFF,
    8'h00, 8'h01, 8'h02, 8'h02, 8'h01, 8'h01, 8'h00, 8'h00,
    8'h00, 8'h02, 8'h03, 8'h00, 8'hFF, 8'hFE, 8'hFE, 8'h00,
    8'h01, 8'h00, 8'h01, 8'h01, 8'hFF, 8'hFF, 8'h02, 8'h00,
    8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00,
    8'h01, 8'h00, 8'h01, 8'h01, 8'hFF, 8'hFF, 8'h00, 8'h00,
    8'hFF, 8'h00, 8'h00, 8'h00, 8'h01, 8'h01, 8'h00, 8'h00,
    8'hFF, 8'hFD, 8'hFE, 8'hFE, 8'hFE, 8'hFD, 8'hFF, 8'hFF,
    8'h00, 8'h00, 8'h00, 8'h00, 8'hFB, 8'hF9, 8'hF9, 8'hFA,
    8'hFB, 8'hFB, 8'hFA, 8'hFB, 8'hFF, 8'hF7, 8'hFE, 8'h01,
    8'hFF, 8'hFF, 8'h00, 8'hFE, 8'hFE, 8'hFE, 8'hFF, 8'hFF,
    8'hFF, 8'h00, 8'hFC, 8'hFB, 8'h04, 8'hFD, 8'h00, 8'hFE,
    8'hFE, 8'hFF, 8'hFE, 8'h01, 8'h01, 8'h00, 8'h01, 8'h00,
    8'hFD, 8'h03, 8'hFF, 8'hFF, 8'hFE, 8'hFE, 8'hFE, 8'h00,
    8'h03, 8'h02, 8'h02, 8'h02, 8'h01, 8'h00, 8'h02, 8'h02,
    8'h00, 8'h00, 8'hFF, 8'hFE, 8'h00, 8'h03, 8'h03, 8'h01,
    8'h01, 8'hFD, 8'hFE, 8'h03, 8'h01, 8'h01, 8'h02, 8'h01,
    8'hFF, 8'hFF, 8'h02, 8'h01, 8'h01, 8'h01, 8'hFE, 8'hFC,
    8'h02, 8'h01, 8'h02, 8'h03, 8'h04, 8'hFE, 8'hFE, 8'hFF,
    8'h02, 8'h01, 8'h02, 8'hFF, 8'hF7, 8'hFE, 8'hFF, 8'h00,
    8'h01, 8'h02, 8'hFE, 8'h00, 8'h00, 8'h02, 8'h02, 8'h00,
    8'hFF, 8'hFF, 8'hFE, 8'h00, 8'hFE, 8'h01, 8'hFF, 8'h01,
    8'h00, 8'h01, 8'h01, 8'h01, 8'hFF, 8'hFC, 8'hFD, 8'hFA,
    8'h00, 8'h00, 8'h01, 8'h02, 8'h01, 8'h01, 8'hFF, 8'h00,
    8'hFF, 8'hFE, 8'hFC, 8'h02, 8'hFB, 8'h01, 8'h03, 8'h02,
    8'h00, 8'h01, 8'h00, 8'h00, 8'hFF, 8'h00, 8'hFF, 8'hFA,
    8'hFF, 8'h01, 8'h02, 8'h00, 8'h01, 8'h02, 8'h00, 8'h02,
    8'h02, 8'h02, 8'h02, 8'h03, 8'h01, 8'hFE, 8'h00, 8'hFF,
    8'hFD, 8'hFA, 8'hFC, 8'hFB, 8'hFB, 8'hFB, 8'hFB, 8'hFD,
    8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'h01, 8'h01, 8'h00,
    8'hFD, 8'hFF, 8'h00, 8'h00, 8'hFC, 8'hF9, 8'hFC, 8'hFC,
    8'h03, 8'hFF, 8'h01, 8'h01, 8'h01, 8'h00, 8'h00, 8'h00,
    8'h02, 8'h00, 8'hFF, 8'hFF, 8'hFB, 8'h02, 8'h01, 8'h01,
    8'h01, 8'h00, 8'h00, 8'h00, 8'h01, 8'h01, 8'h01, 8'h00,
    8'h00, 8'hFF, 8'h01, 8'h01, 8'hFF, 8'hFE, 8'hFF, 8'hFE,
    8'hFF, 8'h00, 8'h01, 8'h00, 8'h01, 8'h00, 8'hFC, 8'h00,
    8'h01, 8'hFF, 8'hFD, 8'hFD, 8'hFA, 8'hFB, 8'hFD, 8'h00,
    8'hFF, 8'h00, 8'hFE, 8'h00, 8'h01, 8'h01, 8'h00, 8'hFC,
    8'hFE, 8'hFE, 8'hFF, 8'hFE, 8'h01, 8'h01, 8'h01, 8'h00,
    8'hFE, 8'h00, 8'h01, 8'hFE, 8'hFE, 8'h01, 8'hFF, 8'hFF,
    8'hFE, 8'h01, 8'h02, 8'h00, 8'hFD, 8'h00, 8'hFF, 8'h00,
    8'h00, 8'h00, 8'h01, 8'hFF, 8'hFF, 8'hFE, 8'hFD, 8'h04,
    8'h00, 8'hFE, 8'h01, 8'hFC, 8'h00, 8'hFE, 8'hFE, 8'hFF,
    8'hFF, 8'hFF, 8'hFD, 8'hFC, 8'hFF, 8'hFD, 8'hFD, 8'hFF,
    8'hF9, 8'hFF, 8'h00, 8'h00, 8'h00, 8'hFF, 8'h00, 8'hFE,
    8'hFC, 8'hFA, 8'hFB, 8'hFC, 8'hFD, 8'hFD, 8'h02, 8'h02,
    8'h00, 8'hFF, 8'hFE, 8'hFE, 8'hFB, 8'hFA, 8'hF9, 8'hFE,
    8'hFC, 8'hFE, 8'h02, 8'hFE, 8'hFF, 8'h02, 8'h04, 8'h03,
    8'h01, 8'h01, 8'h02, 8'h00, 8'h02, 8'h03, 8'h00, 8'h00,
    8'h00, 8'hFE, 8'h00, 8'hFD, 8'hFF, 8'hFE, 8'hFE, 8'hFD,
    8'hFE, 8'hFD, 8'hFE, 8'h00, 8'hFD, 8'hFC, 8'hFB, 8'hFC,
    8'hF9, 8'hFA, 8'hFC, 8'hFC, 8'hFD, 8'h00, 8'hFF, 8'hFF,
    8'hFF, 8'hFD, 8'h04, 8'h04, 8'h03, 8'h02, 8'h04, 8'h04,
    8'h00, 8'h00, 8'hFC, 8'hFD, 8'hFA, 8'hFC, 8'h01, 8'h03,
    8'h03, 8'h03, 8'h04, 8'h02, 8'h01, 8'h01, 8'h00, 8'hFC,
    8'hFC, 8'hFB, 8'hFB, 8'h01, 8'h02, 8'h02, 8'h03, 8'h03,
    8'h01, 8'h02, 8'h01, 8'h00, 8'hFC, 8'hFC, 8'hFD, 8'h00,
    8'h00, 8'h02, 8'h00, 8'h02, 8'h02, 8'h00, 8'h01, 8'hFF,
    8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'h01, 8'h02, 8'h02, 8'hFE,
    8'h00, 8'h02, 8'hFD, 8'hFC, 8'h00, 8'h00, 8'h00, 8'h00,
    8'hFE, 8'h01, 8'h03, 8'hFF, 8'hFE, 8'hFE, 8'h00, 8'hFC,
    8'hFA, 8'hFF, 8'h01, 8'h01, 8'hFE, 8'hFF, 8'hFB, 8'hFD,
    8'hFE, 8'hFD, 8'h00, 8'hFF, 8'hFD, 8'h00, 8'hFF, 8'hFF,
    8'h01, 8'h00, 8'h00, 8'h00, 8'hFE, 8'hFE, 8'hFD, 8'hFE,
    8'hFE, 8'hFD, 8'hFE, 8'hFF, 8'hFF, 8'h00, 8'hFD, 8'hFF,
    8'h03, 8'hF8, 8'hFE, 8'hFD, 8'hFC, 8'hFB, 8'hFC, 8'hFD,
    8'hFE, 8'hFF, 8'hFD, 8'hFF, 8'hFD, 8'hFE, 8'hFB, 8'h00,
    8'hFF, 8'hFC, 8'hFD, 8'hFD, 8'h00, 8'h00, 8'hFE, 8'hFE,
    8'hFD, 8'hFB, 8'h00, 8'h04, 8'h00, 8'h00, 8'h00, 8'hFF,
    8'hFF, 8'h01, 8'h00, 8'h00, 8'h00, 8'hFD, 8'hFB, 8'hFE,
    8'h01, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
    8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
    8'h00, 8'h01, 8'h00, 8'hFF, 8'hFE, 8'hFF, 8'h00, 8'h00,
    8'h01, 8'hFF, 8'h00, 8'hFF, 8'h00, 8'h00, 8'h02, 8'h00,
    8'h00, 8'h00, 8'h00, 8'hFF, 8'h00, 8'h01, 8'h01, 8'h00,
    8'h00, 8'hFE, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'hFE, 8'hFC,
    8'hFE, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF,
    8'hFD, 8'hFC, 8'hFD, 8'hFE, 8'h01, 8'h01, 8'hFE, 8'h00,
    8'h00, 8'h00, 8'h00, 8'hFC, 8'hFA, 8'hF7, 8'hFA, 8'hFA,
    8'hFE, 8'h03, 8'h03, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00,
    8'hFE, 8'hFB, 8'hF8, 8'hF9, 8'hFB, 8'h00, 8'h01, 8'h02,
    8'h01, 8'h01, 8'h00, 8'h00, 8'h01, 8'hFF, 8'hFF, 8'hFD,
    8'hFD, 8'hFD, 8'hFC, 8'hFF, 8'hFE, 8'h00, 8'h00, 8'hFF,
    8'h00, 8'h00, 8'h00, 8'h02, 8'h00, 8'hFE, 8'hFD, 8'hFC,
    8'hFD, 8'hFE, 8'hFD, 8'hFF, 8'h00, 8'h00, 8'h00, 8'hFE,
    8'hFE, 8'hFE, 8'hFA, 8'hFB, 8'hFC, 8'hFD, 8'hFE, 8'hFE,
    8'h00, 8'h00, 8'h00, 8'h00, 8'hFE, 8'hFC, 8'hFD, 8'hFD,
    8'hFE, 8'h00, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h01,
    8'h00, 8'h00, 8'hFE, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00,
    8'h00, 8'hFF, 8'h00, 8'h00, 8'h00, 8'hFF, 8'h00, 8'hFF,
    8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h01,
    8'h00, 8'h00, 8'h00, 8'h00, 8'hFD, 8'hFC, 8'hFE, 8'hFD,
    8'hFC, 8'h00, 8'hFC, 8'hFB, 8'hFF, 8'hFD, 8'hFD, 8'hFE,
    8'hFD, 8'h02, 8'h01, 8'h00, 8'h01, 8'h01, 8'h01, 8'hFE,
    8'h00, 8'hFC, 8'h02, 8'hFD, 8'h00, 8'h01, 8'h02, 8'h01,
    8'h01, 8'h00, 8'h02, 8'h01, 8'h01, 8'hFF, 8'h00, 8'hFF,
    8'hFB, 8'h01, 8'h02, 8'h02, 8'h02, 8'h01, 8'h01, 8'h01,
    8'hFF, 8'h00, 8'hFF, 8'hFF, 8'hFE, 8'h00, 8'h01, 8'h02,
    8'h01, 8'h01, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01,
    8'h01, 8'hFF, 8'hFD, 8'h01, 8'h01, 8'hFF, 8'hFF, 8'hFE,
    8'h00, 8'h00, 8'h01, 8'h02, 8'h02, 8'h03, 8'h02, 8'h02,
    8'hFE, 8'hFF, 8'h00, 8'hFF, 8'h00, 8'h00, 8'h01, 8'h00,
    8'h00, 8'h00, 8'h01, 8'h02, 8'hFC, 8'hFD, 8'h01, 8'h03,
    8'h02, 8'h02, 8'h03, 8'hFF, 8'hFF, 8'hFD, 8'hFC, 8'hFF,
    8'h01, 8'h00, 8'hFF, 8'h02, 8'h02, 8'h04, 8'h03, 8'h01,
    8'hFE, 8'hFD, 8'hFE, 8'hFE, 8'h01, 8'hFC, 8'hF9, 8'hFE,
    8'h00, 8'h01, 8'h02, 8'h02, 8'h01, 8'hFF, 8'h00, 8'h00,
    8'h01, 8'h01, 8'hFB, 8'hFC, 8'hFE, 8'h01, 8'hFF, 8'hFE,
    8'hFF, 8'h00, 8'h01, 8'h00, 8'h01, 8'h01, 8'h01, 8'hFB,
    8'hFC, 8'hFE, 8'hFF, 8'hFD, 8'hFC, 8'hFE, 8'h00, 8'h01,
    8'h01, 8'h01, 8'h02, 8'h02, 8'hFD, 8'hFF, 8'hFE, 8'h00,
    8'hFF, 8'hFE, 8'hFF, 8'hFF, 8'h01, 8'h00, 8'hFD, 8'hFB,
    8'hFB, 8'hFE, 8'h05, 8'h03, 8'h02, 8'h00, 8'h01, 8'hFF,
    8'hFF, 8'hFE, 8'h00, 8'hFE, 8'hFF, 8'h01, 8'hFF, 8'h03,
    8'hFE, 8'h00, 8'h00, 8'hFF, 8'h01, 8'h01, 8'h01, 8'h00,
    8'h00, 8'h00, 8'hFE, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h01,
    8'h01, 8'h01, 8'h01, 8'h02, 8'h02, 8'h02, 8'h01, 8'h02,
    8'hFF, 8'h01, 8'hFF, 8'h01, 8'h01, 8'h01, 8'h02, 8'h02,
    8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h00, 8'hFF, 8'hFF,
    8'h00, 8'h02, 8'h03, 8'h03, 8'h02, 8'h03, 8'h02, 8'h02,
    8'h00, 8'h03, 8'h03, 8'h00, 8'h00, 8'h02, 8'h02, 8'h00,
    8'h03, 8'h00, 8'h02, 8'h02, 8'h01, 8'h02, 8'h00, 8'hFB,
    8'h01, 8'h00, 8'hFE, 8'h01, 8'h03, 8'h03, 8'h01, 8'h02,
    8'h02, 8'h02, 8'h01, 8'hFF, 8'hFD, 8'h00, 8'h01, 8'h00,
    8'h02, 8'h01, 8'h03, 8'h02, 8'h02, 8'h05, 8'hFF, 8'h00,
    8'h00, 8'h01, 8'hFC, 8'hFF, 8'h00, 8'h02, 8'h02, 8'h02,
    8'h00, 8'h02, 8'h02, 8'h00, 8'h01, 8'hFF, 8'hFC, 8'hFD,
    8'hFF, 8'h00, 8'h02, 8'h01, 8'h02, 8'hFF, 8'h01, 8'h00,
    8'h00, 8'h00, 8'h00, 8'hF9, 8'hFD, 8'h00, 8'h00, 8'h02,
    8'h02, 8'h04, 8'h03, 8'h03, 8'h02, 8'h00, 8'h00, 8'hFE,
    8'hFE, 8'hFE, 8'hFF, 8'hFE, 8'hFF, 8'h02, 8'h03, 8'h02,
    8'h04, 8'h01, 8'h02, 8'h00, 8'hFF, 8'hFE, 8'h01, 8'hFF,
    8'hFF, 8'hFD, 8'hFD, 8'hFF, 8'hFE, 8'hFE, 8'hFD, 8'hFC,
    8'hFE, 8'h02, 8'h05, 8'h00, 8'hFE, 8'hFD, 8'hFD, 8'hFC,
    8'h00, 8'hFD, 8'hFF, 8'hFD, 8'hFD, 8'hFE, 8'hFF, 8'h00,
    8'hFC, 8'hFC, 8'hF9, 8'hF9, 8'h00, 8'h02, 8'h02, 8'h01,
    8'h02, 8'h03, 8'h02, 8'h01, 8'h03, 8'hFB, 8'hF6, 8'hFE,
    8'hFE, 8'hFD, 8'h01, 8'h01, 8'h00, 8'h01, 8'h02, 8'h03,
    8'h00, 8'h05, 8'hFE, 8'hFE, 8'hFE, 8'h01, 8'hFE, 8'h01,
    8'h00, 8'h02, 8'h02, 8'h02, 8'h00, 8'h00, 8'hFE, 8'h00,
    8'hFE, 8'hFE, 8'h00, 8'h00, 8'h02, 8'h02, 8'h00, 8'h00,
    8'h01, 8'h02, 8'hFF, 8'h01, 8'hFE, 8'h01, 8'h02, 8'h03,
    8'h01, 8'h02, 8'h02, 8'hFF, 8'hFE, 8'hFF, 8'h00, 8'hFC,
    8'hFF, 8'h01, 8'h00, 8'h02, 8'h01, 8'h01, 8'h01, 8'h01,
    8'h00, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFE, 8'h01,
    8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h01, 8'h03, 8'h01,
    8'h03, 8'h00, 8'hFC, 8'hFE, 8'hFE, 8'hFE, 8'hFC, 8'hFC,
    8'hFF, 8'hFF, 8'h02, 8'h02, 8'h01, 8'hFE, 8'hFC, 8'hFA,
    8'hFE, 8'hFE, 8'hFD, 8'hFC, 8'hFD, 8'h00, 8'h02, 8'h01,
    8'h00, 8'hFE, 8'hFF, 8'h01, 8'hFC, 8'hFE, 8'hFE, 8'hFF,
    8'hFF, 8'hFF, 8'h01, 8'h01, 8'hFF, 8'hFF, 8'hFE, 8'hFE,
    8'hFC, 8'hFB, 8'hFC, 8'hFF, 8'hFF, 8'h00, 8'hFF, 8'h01,
    8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h01, 8'hF9, 8'hFE,
    8'hFE, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'h00, 8'hFF, 8'hFE,
    8'h00, 8'hFF, 8'hFF, 8'hF7, 8'hFF, 8'h00, 8'h00, 8'h00,
    8'hFF, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
    8'h00, 8'hFF, 8'hFF, 8'h00, 8'hFF, 8'h00, 8'h00, 8'h00,
    8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00,
    8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h01, 8'hFF,
    8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h04,
    8'h04, 8'h01, 8'hFE, 8'hFE, 8'hFB, 8'hFD, 8'hFF, 8'h00,
    8'h00, 8'h00, 8'h01, 8'h01, 8'h01, 8'h00, 8'hFF, 8'hFF,
    8'hFE, 8'hFD, 8'hFE, 8'hFE, 8'hFF, 8'h00, 8'hFF, 8'hFE,
    8'hFD, 8'hFC, 8'hFE, 8'hFF, 8'hFD, 8'hFD, 8'hFC, 8'hFC,
    8'hFF, 8'h00, 8'h00, 8'hFD, 8'hFD, 8'hFA, 8'hFB, 8'hFE,
    8'h02, 8'hFD, 8'hFB, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF,
    8'hFE, 8'hFD, 8'hFB, 8'hFC, 8'h02, 8'h03, 8'hFF, 8'hFF,
    8'hFF, 8'h01, 8'h00, 8'hFF, 8'h00, 8'h00, 8'hFE, 8'hFD,
    8'hFE, 8'h03, 8'h02, 8'h01, 8'hFF, 8'hFF, 8'h00, 8'h00,
    8'h00, 8'h00, 8'h00, 8'hFE, 8'h00, 8'h01, 8'h03, 8'h03,
    8'h02, 8'hFF, 8'hFE, 8'h00, 8'h00, 8'hFF, 8'h00, 8'h00,
    8'hFF, 8'h00, 8'h01, 8'h03, 8'h00, 8'hFF, 8'hFF, 8'hFF,
    8'hFF, 8'h00, 8'h00, 8'h00, 8'hFF, 8'h00, 8'h00, 8'hFF,
    8'hFF, 8'hFE, 8'hFD, 8'hFD, 8'hFF, 8'hFF, 8'h00, 8'h00,
    8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF,
    8'hFF, 8'hFE, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00,
    8'hFE, 8'hFF, 8'hFD, 8'hFC, 8'hFA, 8'hFB, 8'hFB, 8'hFC,
    8'hFE, 8'h00, 8'hFF, 8'hFF, 8'hFE, 8'hFB, 8'hF9, 8'h01,
    8'h00, 8'hFF, 8'hFE, 8'hFD, 8'hFF, 8'hF7, 8'hFC, 8'hFF,
    8'hFC, 8'hFA, 8'h01, 8'h02, 8'h02, 8'h01, 8'h00, 8'h00,
    8'hFE, 8'hFF, 8'hFD, 8'hFE, 8'hFC, 8'hFE, 8'h02, 8'h03,
    8'h01, 8'h02, 8'h02, 8'h02, 8'hFF, 8'h00, 8'hFE, 8'hFD,
    8'hFC, 8'hFC, 8'h01, 8'h01, 8'h02, 8'h02, 8'h03, 8'h04,
    8'h02, 8'h01, 8'hFF, 8'hFE, 8'hFD, 8'hFF, 8'hFF, 8'h01,
    8'h01, 8'h02, 8'h01, 8'h01, 8'h01, 8'h02, 8'h01, 8'h01,
    8'h02, 8'h01, 8'hFC, 8'hFE, 8'h03, 8'h00, 8'hFF, 8'hFE,
    8'hFD, 8'h02, 8'h01, 8'h01, 8'h02, 8'h02, 8'h01, 8'hFD,
    8'hFD, 8'h01, 8'hFF, 8'hFD, 8'hFC, 8'hFE, 8'h01, 8'h00,
    8'h00, 8'h03, 8'h01, 8'hFF, 8'hFE, 8'hFF, 8'h00, 8'hFE,
    8'hFD, 8'hFB, 8'hFE, 8'h00, 8'h00, 8'h01, 8'h00, 8'h01,
    8'hFE, 8'hFC, 8'hFE, 8'h00, 8'h01, 8'hFD, 8'hFC, 8'hFD,
    8'hFF, 8'hFF, 8'hFF, 8'h01, 8'hFE, 8'hFF, 8'h01, 8'hF9,
    8'h02, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'h00, 8'h01, 8'hFE,
    8'hFF, 8'h00, 8'hFF, 8'hFD, 8'hFF, 8'h00, 8'h00, 8'h03,
    8'h02, 8'h01, 8'h00, 8'hFF, 8'hFE, 8'h00, 8'h00, 8'h00,
    8'hFE, 8'hFB, 8'h02, 8'h02, 8'h02, 8'h03, 8'h01, 8'h00,
    8'h00, 8'hFF, 8'h02, 8'h00, 8'hFE, 8'h00, 8'h03, 8'h03,
    8'h02, 8'h00, 8'hFD, 8'hFB, 8'hF8, 8'hF6, 8'hFB, 8'h00,
    8'hFE, 8'h02, 8'h04, 8'h03, 8'h02, 8'hFE, 8'hFD, 8'hFF,
    8'h02, 8'h00, 8'hFD, 8'hFE, 8'h01, 8'h00, 8'hF6, 8'hFD,
    8'hFC, 8'hFA, 8'hFE, 8'h00, 8'h01, 8'h01, 8'h02, 8'h03,
    8'h02, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFB, 8'h00, 8'h01,
    8'h00, 8'h02, 8'h03, 8'h04, 8'h04, 8'h01, 8'hFF, 8'h00,
    8'hFE, 8'hFF, 8'h00, 8'h01, 8'h01, 8'h02, 8'h02, 8'h02,
    8'h03, 8'h01, 8'h02, 8'h00, 8'h00, 8'hFE, 8'hFD, 8'h00,
    8'h03, 8'h01, 8'h01, 8'h02, 8'h02, 8'h02, 8'h02, 8'h01,
    8'h00, 8'hFE, 8'hFE, 8'hFC, 8'h00, 8'h00, 8'h00, 8'h00,
    8'h00, 8'hFF, 8'h02, 8'hFF, 8'hFE, 8'hFE, 8'hFC, 8'hF9,
    8'hF5, 8'h00, 8'hFE, 8'h01, 8'h00, 8'h01, 8'h02, 8'h02,
    8'hFE, 8'hFD, 8'hFF, 8'hFC, 8'hFC, 8'hF7, 8'hFE, 8'hFF,
    8'hFD, 8'hFE, 8'h00, 8'h02, 8'h00, 8'hFE, 8'hFE, 8'hFC,
    8'h00, 8'hFE, 8'hFE, 8'hFD, 8'hFE, 8'hFE, 8'h00, 8'h00,
    8'hFF, 8'h01, 8'hFF, 8'hFC, 8'hFC, 8'h00, 8'hFC, 8'h03,
    8'hFE, 8'h02, 8'hFF, 8'h01, 8'h01, 8'h03, 8'h01, 8'hFF,
    8'hFF, 8'hFF, 8'h00, 8'h02, 8'h00, 8'hFF, 8'hFF, 8'h00,
    8'hFE, 8'hFF, 8'h00, 8'hFF, 8'h00, 8'hFE, 8'hFF, 8'hFD,
    8'h03, 8'h02, 8'hFF, 8'h04, 8'h04, 8'h02, 8'h02, 8'h03,
    8'h04, 8'h01, 8'h02, 8'h04, 8'h01, 8'h00, 8'h03, 8'h00,
    8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFC, 8'hFC, 8'hFB,
    8'hFD, 8'hFC, 8'hFF, 8'h01, 8'hFD, 8'hFA, 8'hFD, 8'hFC,
    8'hF9, 8'hF8, 8'hF7, 8'hF9, 8'hFF, 8'hFF, 8'hFB, 8'hFC,
    8'h00, 8'hFB, 8'hFD, 8'hF6, 8'hF3, 8'hFD, 8'h00, 8'h02,
    8'h03, 8'h03, 8'h00, 8'hF8, 8'hF8, 8'hFD, 8'hF8, 8'hF6,
    8'hFA, 8'hFD, 8'hFF, 8'h00, 8'h04, 8'h03, 8'h02, 8'h02,
    8'h03, 8'hFE, 8'hFF, 8'hFF, 8'hFE, 8'hFF, 8'hFD, 8'hFE,
    8'h01, 8'h02, 8'h00, 8'h02, 8'h01, 8'h01, 8'hFF, 8'hF8,
    8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h02, 8'h01, 8'h03, 8'h00,
    8'h03, 8'h00, 8'hFE, 8'h00, 8'hFD, 8'hFF, 8'h00, 8'h01,
    8'h00, 8'h01, 8'h01, 8'h02, 8'h01, 8'hFD, 8'hFE, 8'hFD,
    8'hFF, 8'hFA, 8'hFE, 8'h01, 8'h01, 8'h01, 8'h02, 8'h03,
    8'h00, 8'h01, 8'hFD, 8'hFD, 8'hFF, 8'hFB, 8'hFC, 8'hFC,
    8'h00, 8'h02, 8'h02, 8'h03, 8'h01, 8'hFF, 8'hFF, 8'hFD,
    8'hFB, 8'hFF, 8'hFE, 8'hF8, 8'hFE, 8'hFE, 8'h00, 8'h03,
    8'h03, 8'h00, 8'hFE, 8'hFE, 8'hFD, 8'hFE, 8'hFF, 8'h00,
    8'hFD, 8'hFB, 8'h01, 8'h01, 8'h01, 8'h01, 8'hFF, 8'hFD,
    8'hFD, 8'hFE, 8'h01, 8'h00, 8'h05, 8'h02, 8'hFE, 8'h00,
    8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h00,
    8'h00, 8'h03, 8'hFF, 8'hF9, 8'h03, 8'h00, 8'h00, 8'h01,
    8'h01, 8'h00, 8'h00, 8'h01, 8'h02, 8'h01, 8'h00, 8'hFE
};

