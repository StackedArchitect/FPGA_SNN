// Automatically generated weight parameters for FC_BIAS
// Bit width: 8
// Generated from quantize_weights.py

// Total weights: 10
// Original shape: (10,)

parameter [7:0] FC_BIAS [0:9] = '{
    8'h01, 8'h02, 8'hFF, 8'hFF, 8'h01, 8'hFF, 8'h00, 8'h01,
    8'h00, 8'h00
};

