// Automatically generated weight parameters for CONV_WEIGHTS
// Bit width: 8
// Generated from quantize_weights.py

// Total weights: 36
// Original shape: (4, 1, 3, 3)

parameter [7:0] CONV_WEIGHTS [0:35] = '{
    8'h09, 8'h0B, 8'hFE, 8'h01, 8'hFE, 8'hF5, 8'hEF, 8'hF7,
    8'hF8, 8'hF6, 8'h07, 8'h0A, 8'h00, 8'h0A, 8'hFF, 8'h06,
    8'h04, 8'hF7, 8'hF7, 8'hF2, 8'h06, 8'hFD, 8'hFF, 8'h04,
    8'h0D, 8'h07, 8'hFE, 8'h03, 8'h0A, 8'h09, 8'hF9, 8'h06,
    8'h0B, 8'hF0, 8'hED, 8'hF0
};

